module AsciiToGraph
(
    input [7:0]AC,
    output reg [48:0]col
);
    reg [6:0]C[6:0];
    always@(*)begin
        case(AC)
				8'd0:begin
                C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0000000;
                C[3]=7'b0000000;
                C[4]=7'b0000000;
                C[5]=7'b0000000;
                C[6]=7'b0000000;
            end
				8'd1:begin
                C[0]=7'b1111111;
                C[1]=7'b1111111;
                C[2]=7'b1111111;
                C[3]=7'b1111111;
                C[4]=7'b1111111;
                C[5]=7'b1111111;
                C[6]=7'b1111111;
            end
            8'd48:begin
                C[0]=7'b0011100;
                C[1]=7'b0100010;
                C[2]=7'b0100110;
                C[3]=7'b0101010;
                C[4]=7'b0110010;
                C[5]=7'b0100010;
                C[6]=7'b0011100;
            end
            8'd49:begin
                C[0]=7'b0001000;
                C[1]=7'b0011000;
                C[2]=7'b0001000;
                C[3]=7'b0001000;
                C[4]=7'b0001000;
                C[5]=7'b0001000;
                C[6]=7'b0011100;
            end
				8'd50:begin
			       C[0]=7'b0011100;
                C[1]=7'b0100010;
                C[2]=7'b0000010;
                C[3]=7'b0000100;
                C[4]=7'b0001000;
                C[5]=7'b0010000;
                C[6]=7'b0111110;
				end
				8'd51:begin
					 C[0]=7'b0111110;
                C[1]=7'b0000100;
                C[2]=7'b0001000;
                C[3]=7'b0000100;
                C[4]=7'b0000010;
                C[5]=7'b0100010;
                C[6]=7'b0011100;
				end
				8'd52:begin
					 C[0]=7'b0000100;
                C[1]=7'b0001100;
                C[2]=7'b0010100;
                C[3]=7'b0100100;
                C[4]=7'b0111110;
                C[5]=7'b0000100;
                C[6]=7'b0000100;
				end
				8'd53:begin
					 C[0]=7'b0111110;
                C[1]=7'b0100000;
                C[2]=7'b0111100;
                C[3]=7'b0000010;
                C[4]=7'b0000010;
                C[5]=7'b0100010;
                C[6]=7'b0011100;
				end
				8'd54:begin
					 C[0]=7'b0001100;
                C[1]=7'b0010000;
                C[2]=7'b0100000;
                C[3]=7'b0111100;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0011100;
				end
				8'd55:begin
					 C[0]=7'b0111110;
                C[1]=7'b0000010;
                C[2]=7'b0000100;
                C[3]=7'b0001000;
                C[4]=7'b0010000;
                C[5]=7'b0010000;
                C[6]=7'b0010000;
				end
				8'd56:begin
					 C[0]=7'b0011100;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0011100;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0011100;					 
				end
				8'd57:begin
				    C[0]=7'b0011100;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0011110;
                C[4]=7'b0000010;
                C[5]=7'b0000100;
                C[6]=7'b0011000;
				end
				8'd65:begin
				    C[0]=7'b0011100;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0100010;
                C[4]=7'b0111110;
                C[5]=7'b0100010;
                C[6]=7'b0100010;
				end
				8'd66:begin
				    C[0]=7'b0111100;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0111100;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0111100;
				end
				8'd67:begin
				    C[0]=7'b0011100;
                C[1]=7'b0100010;
                C[2]=7'b0100000;
                C[3]=7'b0100000;
                C[4]=7'b0100000;
                C[5]=7'b0100010;
                C[6]=7'b0011100;
				end
				8'd68:begin
				    C[0]=7'b0111000;
                C[1]=7'b0100100;
                C[2]=7'b0100010;
                C[3]=7'b0100010;
                C[4]=7'b0100010;
                C[5]=7'b0100100;
                C[6]=7'b0111000;
				end
				8'd69:begin
				    C[0]=7'b0111110;
                C[1]=7'b0100000;
                C[2]=7'b0100000;
                C[3]=7'b0111100;
                C[4]=7'b0100000;
                C[5]=7'b0100000;
                C[6]=7'b0111110;
				end
				8'd70:begin
				    C[0]=7'b0111110;
                C[1]=7'b0100000;
                C[2]=7'b0100000;
                C[3]=7'b0111100;
                C[4]=7'b0100000;
                C[5]=7'b0100000;
                C[6]=7'b0100000;
				end
				8'd71:begin
				    C[0]=7'b0011100;
                C[1]=7'b0100010;
                C[2]=7'b0100000;
                C[3]=7'b0101110;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0011110;
				end
				8'd72:begin
				    C[0]=7'b0100010;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0111110;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0100010;
				end
				8'd73:begin
				    C[0]=7'b0011100;
                C[1]=7'b0001000;
                C[2]=7'b0001000;
                C[3]=7'b0001000;
                C[4]=7'b0001000;
                C[5]=7'b0001000;
                C[6]=7'b0011100;
				end
				8'd74:begin
				    C[0]=7'b0001110;
                C[1]=7'b0000100;
                C[2]=7'b0000100;
                C[3]=7'b0000100;
                C[4]=7'b0000100;
                C[5]=7'b0100100;
                C[6]=7'b0011000;
				end
				8'd75:begin
				    C[0]=7'b0100010;
                C[1]=7'b0100100;
                C[2]=7'b0101000;
                C[3]=7'b0110000;
                C[4]=7'b0101000;
                C[5]=7'b0100100;
                C[6]=7'b0100010;
				end
				8'd76:begin
				    C[0]=7'b0100000;
                C[1]=7'b0100000;
                C[2]=7'b0100000;
                C[3]=7'b0100000;
                C[4]=7'b0100000;
                C[5]=7'b0100000;
                C[6]=7'b0111110;
				end
				8'd77:begin
				    C[0]=7'b0100010;
                C[1]=7'b0110110;
                C[2]=7'b0101010;
                C[3]=7'b0101010;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0100010;
				end
				8'd78:begin
				    C[0]=7'b0100010;
                C[1]=7'b0100010;
                C[2]=7'b0110010;
                C[3]=7'b0101010;
                C[4]=7'b0100110;
                C[5]=7'b0100010;
                C[6]=7'b0100010;
				end
				8'd79:begin
				    C[0]=7'b0011100;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0100010;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0011100;
				end
				8'd80:begin
				    C[0]=7'b0111100;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0111100;
                C[4]=7'b0100000;
                C[5]=7'b0100000;
                C[6]=7'b0100000;
				end
				8'd81:begin
				    C[0]=7'b0011100;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0100010;
                C[4]=7'b0101010;
                C[5]=7'b0100100;
                C[6]=7'b0011010;
				end
				8'd82:begin
				    C[0]=7'b0111100;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0111100;
                C[4]=7'b0101000;
                C[5]=7'b0100100;
                C[6]=7'b0100010;
				end
				8'd83:begin
				    C[0]=7'b0011110;
                C[1]=7'b0100000;
                C[2]=7'b0100000;
                C[3]=7'b0011100;
                C[4]=7'b0000010;
                C[5]=7'b0000010;
                C[6]=7'b0111100;
				end
				8'd84:begin
				    C[0]=7'b0111110;
                C[1]=7'b0001000;
                C[2]=7'b0001000;
                C[3]=7'b0001000;
                C[4]=7'b0001000;
                C[5]=7'b0001000;
                C[6]=7'b0001000;
				end
				8'd85:begin
				    C[0]=7'b0100010;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0100010;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0011100;
				end
				8'd86:begin
				    C[0]=7'b0100010;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0100010;
                C[4]=7'b0100010;
                C[5]=7'b0010100;
                C[6]=7'b0001000;
				end
				8'd87:begin
				    C[0]=7'b0100010;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0101010;
                C[4]=7'b0101010;
                C[5]=7'b0101010;
                C[6]=7'b0010100;
				end
				8'd88:begin
				    C[0]=7'b0100010;
                C[1]=7'b0100010;
                C[2]=7'b0010100;
                C[3]=7'b0001000;
                C[4]=7'b0010100;
                C[5]=7'b0100010;
                C[6]=7'b0100010;
				end
				8'd89:begin
				    C[0]=7'b0100010;
                C[1]=7'b0100010;
                C[2]=7'b0100010;
                C[3]=7'b0010100;
                C[4]=7'b0001000;
                C[5]=7'b0001000;
                C[6]=7'b0001000;
				end
				8'd90:begin
				    C[0]=7'b0111110;
                C[1]=7'b0000010;
                C[2]=7'b0000100;
                C[3]=7'b0001000;
                C[4]=7'b0010000;
                C[5]=7'b0100000;
                C[6]=7'b0111110;
				end
				8'd33:begin
				    C[0]=7'b0001000;
                C[1]=7'b0001000;
                C[2]=7'b0001000;
                C[3]=7'b0001000;
                C[4]=7'b0001000;
                C[5]=7'b0000000;
                C[6]=7'b0001000;
				end
				8'd34:begin
				    C[0]=7'b0010100;
                C[1]=7'b0010100;
                C[2]=7'b0010100;
                C[3]=7'b0000000;
                C[4]=7'b0000000;
                C[5]=7'b0000000;
                C[6]=7'b0000000;
				end
				8'd35:begin
				    C[0]=7'b0010100;
                C[1]=7'b0010100;
                C[2]=7'b0111110;
                C[3]=7'b0010100;
                C[4]=7'b0111110;
                C[5]=7'b0010100;
                C[6]=7'b0010100;
				end
				8'd36:begin
				    C[0]=7'b0001000;
                C[1]=7'b0011110;
                C[2]=7'b0101000;
                C[3]=7'b0011100;
                C[4]=7'b0001010;
                C[5]=7'b0111100;
                C[6]=7'b0001000;
				end
				8'd37:begin
				    C[0]=7'b0110000;
                C[1]=7'b0110010;
                C[2]=7'b0000100;
                C[3]=7'b0001000;
                C[4]=7'b0010000;
                C[5]=7'b0100110;
                C[6]=7'b0000110;
				end
				8'd38:begin
				    C[0]=7'b0011000;
                C[1]=7'b0100100;
                C[2]=7'b0101000;
                C[3]=7'b0010000;
                C[4]=7'b0101010;
                C[5]=7'b0100100;
                C[6]=7'b0011010;
				end
				8'd39:begin
				    C[0]=7'b0011000;
                C[1]=7'b0001000;
                C[2]=7'b0010000;
                C[3]=7'b0000000;
                C[4]=7'b0000000;
                C[5]=7'b0000000;
                C[6]=7'b0000000;
				end
				8'd40:begin
				    C[0]=7'b0000100;
                C[1]=7'b0001000;
                C[2]=7'b0010000;
                C[3]=7'b0010000;
                C[4]=7'b0010000;
                C[5]=7'b0001000;
                C[6]=7'b0000100;
				end
				8'd41:begin
				    C[0]=7'b0010000;
                C[1]=7'b0001000;
                C[2]=7'b0000100;
                C[3]=7'b0000100;
                C[4]=7'b0000100;
                C[5]=7'b0001000;
                C[6]=7'b0010000;
				end
				8'd42:begin
				    C[0]=7'b0000000;
                C[1]=7'b0001000;
                C[2]=7'b0101010;
                C[3]=7'b0011100;
                C[4]=7'b0101010;
                C[5]=7'b0001000;
                C[6]=7'b0000000;
				end
				8'd43:begin
				    C[0]=7'b0000000;
                C[1]=7'b0001000;
                C[2]=7'b0001000;
                C[3]=7'b0111110;
                C[4]=7'b0001000;
                C[5]=7'b0001000;
                C[6]=7'b0000000;
				end
				8'd44:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0000000;
                C[3]=7'b0000000;
                C[4]=7'b0011000;
                C[5]=7'b0001000;
                C[6]=7'b0010000;
				end
				8'd45:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0000000;
                C[3]=7'b0111110;
                C[4]=7'b0000000;
                C[5]=7'b0000000;
                C[6]=7'b0000000;
				end
				8'd46:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0000000;
                C[3]=7'b0000000;
                C[4]=7'b0000000;
                C[5]=7'b0110000;
                C[6]=7'b0110000;
				end
				8'd47:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000010;
                C[2]=7'b0000100;
                C[3]=7'b0001000;
                C[4]=7'b0010000;
                C[5]=7'b0100000;
                C[6]=7'b0000000;
				end
				8'd58:begin
				    C[0]=7'b0000000;
                C[1]=7'b0011000;
                C[2]=7'b0011000;
                C[3]=7'b0000000;
                C[4]=7'b0011000;
                C[5]=7'b0011000;
                C[6]=7'b0000000;
				end
				8'd59:begin
				    C[0]=7'b0000000;
                C[1]=7'b0011000;
                C[2]=7'b0011000;
                C[3]=7'b0000000;
                C[4]=7'b0011000;
                C[5]=7'b0001000;
                C[6]=7'b0010000;
				end
				8'd60:begin
				    C[0]=7'b0000100;
                C[1]=7'b0001000;
                C[2]=7'b0010000;
                C[3]=7'b0100000;
                C[4]=7'b0010000;
                C[5]=7'b0001000;
                C[6]=7'b0000100;
				end
				8'd61:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0111110;
                C[3]=7'b0000000;
                C[4]=7'b0111110;
                C[5]=7'b0000000;
                C[6]=7'b0000000;
				end
				8'd62:begin
				    C[0]=7'b0010000;
                C[1]=7'b0001000;
                C[2]=7'b0000100;
                C[3]=7'b0000010;
                C[4]=7'b0000100;
                C[5]=7'b0001000;
                C[6]=7'b0010000;
				end
				8'd58:begin
				    C[0]=7'b0011100;
                C[1]=7'b0100010;
                C[2]=7'b0000010;
                C[3]=7'b0000100;
                C[4]=7'b0001000;
                C[5]=7'b0000000;
                C[6]=7'b0001000;
				end
				8'd91:begin
				    C[0]=7'b0111000;
                C[1]=7'b0100000;
                C[2]=7'b0100000;
                C[3]=7'b0100000;
                C[4]=7'b0100000;
                C[5]=7'b0100000;
                C[6]=7'b0111000;
				end
				8'd92:begin
				    C[0]=7'b0100010;
                C[1]=7'b0010100;
                C[2]=7'b0111110;
                C[3]=7'b0001000;
                C[4]=7'b0111110;
                C[5]=7'b0001000;
                C[6]=7'b0001000;
				end
				8'd93:begin
				    C[0]=7'b0011100;
                C[1]=7'b0000100;
                C[2]=7'b0000100;
                C[3]=7'b0000100;
                C[4]=7'b0000100;
                C[5]=7'b0000100;
                C[6]=7'b0011100;
				end
				8'd94:begin
				    C[0]=7'b0001000;
                C[1]=7'b0010100;
                C[2]=7'b0100010;
                C[3]=7'b0000000;
                C[4]=7'b0000000;
                C[5]=7'b0000000;
                C[6]=7'b0000000;
				end
				8'd95:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0000000;
                C[3]=7'b0000000;
                C[4]=7'b0000000;
                C[5]=7'b0000000;
                C[6]=7'b0111110;
				end
				8'd96:begin
				    C[0]=7'b0010000;
                C[1]=7'b0001000;
                C[2]=7'b0000100;
                C[3]=7'b0000000;
                C[4]=7'b0000000;
                C[5]=7'b0000000;
                C[6]=7'b0000000;
				end
				8'd123:begin
				    C[0]=7'b0000100;
                C[1]=7'b0001000;
                C[2]=7'b0001000;
                C[3]=7'b0010000;
                C[4]=7'b0001000;
                C[5]=7'b0001000;
                C[6]=7'b0000100;
				end
				8'd124:begin
				    C[0]=7'b0001000;
                C[1]=7'b0001000;
                C[2]=7'b0001000;
                C[3]=7'b0001000;
                C[4]=7'b0001000;
                C[5]=7'b0001000;
                C[6]=7'b0001000;
				end
				8'd125:begin
				    C[0]=7'b0000000;
                C[1]=7'b0001000;
                C[2]=7'b0000100;
                C[3]=7'b0111110;
                C[4]=7'b0000100;
                C[5]=7'b0001000;
                C[6]=7'b0000000;
				end
				8'd126:begin
				    C[0]=7'b0000000;
                C[1]=7'b0001000;
                C[2]=7'b0010000;
                C[3]=7'b0111110;
                C[4]=7'b0010000;
                C[5]=7'b0001000;
                C[6]=7'b0000000;
				end
				//小寫英文
				8'd97:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0011100;
                C[3]=7'b0000010;
                C[4]=7'b0011110;
                C[5]=7'b0100010;
                C[6]=7'b0011110;
				end
				8'd98:begin
				    C[0]=7'b0100000;
                C[1]=7'b0100000;
                C[2]=7'b0101100;
                C[3]=7'b0110010;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0111100;
				end
				8'd99:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0011100;
                C[3]=7'b0100000;
                C[4]=7'b0100000;
                C[5]=7'b0100010;
                C[6]=7'b0011100;
				end
				8'd100:begin
				    C[0]=7'b0000010;
                C[1]=7'b0000010;
                C[2]=7'b0011010;
                C[3]=7'b0100110;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0011110;
				end
				8'd101:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0011100;
                C[3]=7'b0100010;
                C[4]=7'b0111110;
                C[5]=7'b0100000;
                C[6]=7'b0011100;
				end
				8'd102:begin
				    C[0]=7'b0001100;
                C[1]=7'b0010010;
                C[2]=7'b0010000;
                C[3]=7'b0111000;
                C[4]=7'b0010000;
                C[5]=7'b0010000;
                C[6]=7'b0010000;
				end
				8'd103:begin
				    C[0]=7'b0000000;
                C[1]=7'b0011110;
                C[2]=7'b0100010;
                C[3]=7'b0100010;
                C[4]=7'b0011110;
                C[5]=7'b0000010;
                C[6]=7'b0011100;
				end
				8'd104:begin
				    C[0]=7'b0100000;
                C[1]=7'b0100000;
                C[2]=7'b0101100;
                C[3]=7'b0110010;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0100010;
				end
				8'd105:begin
				    C[0]=7'b0001000;
                C[1]=7'b0000000;
                C[2]=7'b0011000;
                C[3]=7'b0001000;
                C[4]=7'b0001000;
                C[5]=7'b0001000;
                C[6]=7'b0011100;
				end
				8'd106:begin
				    C[0]=7'b0000100;
                C[1]=7'b0000000;
                C[2]=7'b0001100;
                C[3]=7'b0000100;
                C[4]=7'b0000100;
                C[5]=7'b0100100;
                C[6]=7'b0011000;
				end
				8'd107:begin
				    C[0]=7'b0100000;
                C[1]=7'b0100000;
                C[2]=7'b0100100;
                C[3]=7'b0101000;
                C[4]=7'b0110000;
                C[5]=7'b0101000;
                C[6]=7'b0100100;
				end
				8'd108:begin
				    C[0]=7'b0011000;
                C[1]=7'b0001000;
                C[2]=7'b0001000;
                C[3]=7'b0001000;
                C[4]=7'b0001000;
                C[5]=7'b0001000;
                C[6]=7'b0011100;
				end
				8'd109:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0110100;
                C[3]=7'b0101010;
                C[4]=7'b0101010;
                C[5]=7'b0100010;
                C[6]=7'b0100010;
				end
				8'd110:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0101100;
                C[3]=7'b0110010;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0100010;
				end
				8'd111:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0011100;
                C[3]=7'b0100010;
                C[4]=7'b0100010;
                C[5]=7'b0100010;
                C[6]=7'b0011100;
				end
				8'd112:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0111100;
                C[3]=7'b0100010;
                C[4]=7'b0111100;
                C[5]=7'b0100000;
                C[6]=7'b0100000;
				end
				8'd113:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0011010;
                C[3]=7'b0100110;
                C[4]=7'b001110;
                C[5]=7'b0000010;
                C[6]=7'b0000010;
				end
				8'd114:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0101100;
                C[3]=7'b0110010;
                C[4]=7'b0100000;
                C[5]=7'b0100000;
                C[6]=7'b0100000;
				end
				8'd115:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0011100;
                C[3]=7'b0100000;
                C[4]=7'b0011100;
                C[5]=7'b0000010;
                C[6]=7'b0111100;
				end
				8'd116:begin
				    C[0]=7'b0010000;
                C[1]=7'b0010000;
                C[2]=7'b0111000;
                C[3]=7'b0010000;
                C[4]=7'b0010000;
                C[5]=7'b0010010;
                C[6]=7'b0001100;
				end
				8'd117:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0100010;
                C[3]=7'b0100010;
                C[4]=7'b0100010;
                C[5]=7'b0100110;
                C[6]=7'b0011010;
				end
				8'd118:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0100010;
                C[3]=7'b0100010;
                C[4]=7'b0100010;
                C[5]=7'b0010100;
                C[6]=7'b0001000;
				end
				8'd119:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0100010;
                C[3]=7'b0100010;
                C[4]=7'b0101010;
                C[5]=7'b0101010;
                C[6]=7'b0010100;
				end
				8'd120:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0100010;
                C[3]=7'b0010100;
                C[4]=7'b0001000;
                C[5]=7'b0010100;
                C[6]=7'b0100010;
				end
				8'd130:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0100010;
                C[3]=7'b0100010;
                C[4]=7'b0011110;
                C[5]=7'b0000010;
                C[6]=7'b0011100;
				end
				8'd58:begin
				    C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0111110;
                C[3]=7'b0000100;
                C[4]=7'b0001000;
                C[5]=7'b0010000;
                C[6]=7'b0111110;
				end
				default:begin
					 C[0]=7'b0000000;
                C[1]=7'b0000000;
                C[2]=7'b0000000;
                C[3]=7'b0000000;
                C[4]=7'b0000000;
                C[5]=7'b0000000;
                C[6]=7'b0000000;
				end
			endcase
			col={C[0],C[1],C[2],C[3],C[4],C[5],C[6]};
		end
endmodule